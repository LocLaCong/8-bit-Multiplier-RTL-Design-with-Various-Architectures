module WAlLACE (input[7:0] A, input[7:0] B,output[15:0] P);

    reg[7:0] X[7:0];
    integer i, j;
    
reg [7:0]a,b;
initial begin
a=200;b=190;
#10 a=144;b=89;
#10 a=20;b=50;
#10 a=249;b=153;
#10 a=80;b=255;
#10 a=189;b=190;
#10 a=255;b=255;
#10 a=2;b=223;
end
assign A=a,B=b;
   
    always @(A, B) begin
        for(i = 0;i < 8;i = i+1)
            for(j = 0;j < 8;j = j+1)
                X[i][j] <= A[i] & B[j];
    end
    
    wire [52:0]s,c;
    
//redution 8 sang 6

//nhom I

HA HA_0(c[0], s[0], X[0][1], X[1][0]);
FA FA_1(c[1], s[1], X[0][2], X[1][1], X[2][0]);
FA FA_2(c[2], s[2], X[0][3], X[1][2], X[2][1]);
FA FA_3(c[3], s[3], X[0][4], X[1][3], X[2][2]);
FA FA_4(c[4], s[4], X[0][5], X[1][4], X[2][3]);
FA FA_5(c[5], s[5], X[0][6], X[1][5], X[2][4]);
FA FA_6(c[6], s[6], X[0][7], X[1][6], X[2][5]);
HA HA_7(c[7], s[7], X[1][7], X[2][6]);

//nhom II

HA HA_8(c[8], s[8], X[3][1], X[4][0]);
FA FA_9(c[9], s[9], X[3][2], X[4][1], X[5][0]);
FA FA_10(c[10], s[10], X[3][3], X[4][2], X[5][1]);
FA FA_11(c[11], s[11], X[3][4], X[4][3], X[5][2]);
FA FA_12(c[12], s[12], X[3][5], X[4][4], X[5][3]);
FA FA_13(c[13], s[13], X[3][6], X[4][5], X[5][4]);
FA FA_14(c[14], s[14], X[3][7], X[4][6], X[5][5]);
HA HA_15(c[15], s[15], X[4][7], X[5][6]);

//reduction 6 sang 4

//nhom III

HA HA_16(c[16], s[16], s[1], c[0]);
FA FA_17(c[17], s[17], s[2], c[1], X[3][0]);
FA FA_18(c[18], s[18], s[3], c[2], s[8]);
FA FA_19(c[19], s[19], s[4], c[3], s[9]);
FA FA_20(c[20], s[20], s[5], c[4], s[10]);
FA FA_21(c[21], s[21], s[6], c[5], s[11]);
FA FA_22(c[22], s[22], s[7], c[6], s[12]);
FA FA_23(c[23], s[23], X[2][7], c[7], s[13]);

//mhom IV

HA HA_24(c[24], s[24], c[9], X[6][0]);
FA FA_25(c[25], s[25], c[10], X[6][1], X[7][0]);
FA FA_26(c[26], s[26], c[11], X[6][2], X[7][1]);
FA FA_27(c[27], s[27], c[12], X[6][3], X[7][2]);
FA FA_28(c[28], s[28], c[13], X[6][4], X[7][3]);
FA FA_29(c[29], s[29], c[14], X[6][5], X[7][4]);
FA FA_30(c[30], s[30], c[15], X[6][6], X[7][5]);
HA HA_31(c[31], s[31], X[6][7], X[7][6]);

//redution 4 sang 3

//nhom V

HA HA_32(c[32], s[32], s[17], c[16]);
HA HA_33(c[33], s[33], s[18], c[17]);
FA FA_34(c[34], s[34], s[19], c[18], c[8]);
FA FA_35(c[35], s[35], s[20], c[19], s[24]);
FA FA_36(c[36], s[36], s[21], c[20], s[25]);
FA FA_37(c[37], s[37], s[22], c[21], s[26]);
FA FA_38(c[38], s[38], s[23], c[22], s[27]);
FA FA_39(c[39], s[39], s[14], c[23], s[28]);
HA HA_40(c[40], s[40], s[15], s[29]);
HA HA_41(c[41], s[41], X[5][7], s[30]);

//reduction 3 sang 2

//nhom VI

HA HA_42(c[42], s[42], s[33], c[32]);
HA HA_43(c[43], s[43], s[34], c[33]);
HA HA_44(c[44], s[44], s[35], c[34]);
FA FA_45(c[45], s[45], s[36], c[35], c[24]);
FA FA_46(c[46], s[46], s[37], c[36], c[25]);
FA FA_47(c[47], s[47], s[38], c[37], c[26]);
FA FA_48(c[48], s[48], s[39], c[38], c[27]);
FA FA_49(c[49], s[49], s[40], c[39], c[28]);
FA FA_50(c[50], s[50], s[41], c[40], c[29]);
FA FA_51(c[51], s[51], s[31], c[41], c[30]);
HA HA_52(c[52], s[52], X[7][7], c[31]);

//dung bo cong CLA de cong hai so cuoi

wire [10:0]l;
CLA  L10({1'b0,s[52:43]},c[52:42],l); 


assign P = {l,s[42],s[32],s[16],s[0],X[0][0]};

endmodule