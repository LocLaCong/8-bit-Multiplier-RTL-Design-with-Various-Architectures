module CLA(input [10:0]A,B,output[10:0]S);
wire [10:0]G,P;
//Tinh Generate
and Gate1(G[0],A[0],B[0]),
    Gate2(G[1],A[1],B[1]),
    Gate3(G[2],A[2],B[2]),
    Gate4(G[3],A[3],B[3]),
    Gate5(G[4],A[4],B[4]),
    Gate6(G[5],A[5],B[5]),
    Gate7(G[6],A[6],B[6]),
    Gate8(G[7],A[7],B[7]),
    Gate9(G[8],A[8],B[8]),
    Gate10(G[9],A[9],B[9]),
    Gate11(G[10],A[10],B[10]);
//Tinh Propagate
xor Gate12 (P[0],A[0],B[0]),
    Gate13(P[1],A[1],B[1]),
    Gate14(P[2],A[2],B[2]),
    Gate15(P[3],A[3],B[3]),
    Gate16(P[4],A[4],B[4]),
    Gate17(P[5],A[5],B[5]),
    Gate18(P[6],A[6],B[6]),
    Gate19(P[7],A[7],B[7]),
    Gate20(P[8],A[8],B[8]),
    Gate21(P[9],A[9],B[9]),
    Gate22(P[10],A[10],B[10]);
wire [9:0]C;
//Tinh Cout	
assign 
C[0]=G[0], 					
C[1]=G[1]|(P[1]&G[0]),			
C[2]=G[2]|(P[2]&G[1])|(P[2]&P[1]&G[0]),
C[3]=G[3]|(P[3]&G[2])|(P[3]&P[2]&G[1])|(P[3]&P[2]&P[1]&G[0]),
C[4]=G[4]|(P[4]&G[3])|(P[4]&P[3]&G[2])|(P[4]&P[3]&P[2]&G[1])|(P[4]&P[3]&P[2]&P[1]&G[0]),
C[5]=G[5]|(P[5]&G[4])|(P[5]&P[4]&G[3])|(P[5]&P[4]&P[3]&G[2])|(P[5]&P[4]&P[3]&P[2]&G[1])|(P[5]&P[4]&P[3]&P[2]&P[1]&G[0]),
C[6]=G[6]|(P[6]&G[5])|(P[6]&P[5]&G[4])|(P[6]&P[5]&P[4]&G[3])|(P[6]&P[5]&P[4]&P[3]&G[2])|(P[6]&P[5]&P[4]&P[3]&P[2]&G[1])|(P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]),
C[7]=G[7]|(P[7]&G[6])|(P[7]&P[6]&G[5])|(P[7]&P[6]&P[5]&G[4])|(P[7]&P[6]&P[5]&P[4]&G[3])|(P[7]&P[6]&P[5]&P[4]&P[3]&G[2])|(P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1])|(P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]),
C[8]=G[8]|(P[8]&G[7])|(P[8]&P[7]&G[6])|(P[8]&P[7]&P[6]&G[5])|(P[8]&P[7]&P[6]&P[5]&G[4])|(P[8]&P[7]&P[6]&P[5]&P[4]&G[3])|(P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2])|(P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1])|(P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]),
C[9]=G[9]|(P[9]&G[8])|(P[9]&P[8]&G[7])|(P[9]&P[8]&P[7]&G[6])|(P[9]&P[8]&P[7]&P[6]&G[5])|(P[9]&P[8]&P[7]&P[6]&P[5]&G[4])|(P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3])|(P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2])|(P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1])|(P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]);
//C[10]=G[10]|(P[10]&G[9])|(P[10]&P[9]&G[8])|(P[10]&P[9]&P[8]&G[7])|(P[10]&P[9]&P[8]&P[7]&G[6])|(P[10]&P[9]&P[8]&P[7]&P[6]&G[5])|(P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4])|(P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3])|(P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2])|(P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1])|(P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]);

//Tinh S[i]=P[i]^C[i-1];
assign 
S[0]=P[0],
S[1]=P[1]^C[0],
S[2]=P[2]^C[1],
S[3]=P[3]^C[2],
S[4]=P[4]^C[3],
S[5]=P[5]^C[4],
S[6]=P[6]^C[5],
S[7]=P[7]^C[6],
S[8]=P[8]^C[7],
S[9]=P[9]^C[8],
S[10]=P[10]^C[9];
endmodule