module CLA_8bit(input [7:0]A,B,output[8:0]S);
wire [7:0]G,P;

/*reg [7:0]a,b;
initial begin
a=200;b=190;
#10 a=144;b=89;
#10 a=20;b=50;
#10 a=249;b=153;
#10 a=80;b=255;
#10 a=189;b=190;
#10 a=255;b=255;
#10 a=2;b=223;
end
assign A=a,B=b;*/

//G
assign
    G[0]=A[0]&B[0],
    G[1]=A[1]&B[1],
    G[2]=A[2]&B[2],
    G[3]=A[3]&B[3],
    G[4]=A[4]&B[4],
    G[5]=A[5]&B[5],
    G[6]=A[6]&B[6],
    G[7]=A[7]&B[7];
//P
assign
    P[0]=A[0]^B[0],
    P[1]=A[1]^B[1],
    P[2]=A[2]^B[2],
    P[3]=A[3]^B[3],
    P[4]=A[4]^B[4],
    P[5]=A[5]^B[5],
    P[6]=A[6]^B[6],
    P[7]=A[7]^B[7];
wire [7:0]C;

//C[i]=G[i]+P[i]*C[i-1]
assign 
C[0]=G[0], 					
C[1]=G[1]|(P[1]&G[0]),			
C[2]=G[2]|(P[2]&G[1])|(P[2]&P[1]&G[0]),
C[3]=G[3]|(P[3]&G[2])|(P[3]&P[2]&G[1])|(P[3]&P[2]&P[1]&G[0]),
C[4]=G[4]|(P[4]&G[3])|(P[4]&P[3]&G[2])|(P[4]&P[3]&P[2]&G[1])|(P[4]&P[3]&P[2]&P[1]&G[0]),
C[5]=G[5]|(P[5]&G[4])|(P[5]&P[4]&G[3])|(P[5]&P[4]&P[3]&G[2])|(P[5]&P[4]&P[3]&P[2]&G[1])|(P[5]&P[4]&P[3]&P[2]&P[1]&G[0]),
C[6]=G[6]|(P[6]&G[5])|(P[6]&P[5]&G[4])|(P[6]&P[5]&P[4]&G[3])|(P[6]&P[5]&P[4]&P[3]&G[2])|(P[6]&P[5]&P[4]&P[3]&P[2]&G[1])|(P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]),
C[7]=G[7]|(P[7]&G[6])|(P[7]&P[6]&G[5])|(P[7]&P[6]&P[5]&G[4])|(P[7]&P[6]&P[5]&P[4]&G[3])|(P[7]&P[6]&P[5]&P[4]&P[3]&G[2])|(P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1])|(P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]);

//S[i]=P[i]^C[i-1];
assign 
S[0]=P[0],
S[1]=P[1]^C[0],
S[2]=P[2]^C[1],
S[3]=P[3]^C[2],
S[4]=P[4]^C[3],
S[5]=P[5]^C[4],
S[6]=P[6]^C[5],
S[7]=P[7]^C[6],
S[8]=C[7];
endmodule
